module Image_Generator (
    input  i_clk,
    input  i_rst_n
);
endmodule