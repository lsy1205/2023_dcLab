// AltPLL.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module AltPLL (
		output wire  altpll_100k_clk, // altpll_100k.clk
		output wire  altpll_12m_clk,  //  altpll_12m.clk
		output wire  altpll_50m_clk,  //  altpll_50m.clk
		output wire  altpll_800k_clk, // altpll_800k.clk
		input  wire  i_clk_clk,       //       i_clk.clk
		input  wire  i_reset_reset    //     i_reset.reset
	);

	AltPLL_altpll_0 altpll_0 (
		.clk       (i_clk_clk),       //       inclk_interface.clk
		.reset     (i_reset_reset),   // inclk_interface_reset.reset
		.read      (),                //             pll_slave.read
		.write     (),                //                      .write
		.address   (),                //                      .address
		.readdata  (),                //                      .readdata
		.writedata (),                //                      .writedata
		.c0        (altpll_50m_clk),  //                    c0.clk
		.c1        (altpll_12m_clk),  //                    c1.clk
		.c2        (altpll_100k_clk), //                    c2.clk
		.c3        (altpll_800k_clk), //                    c3.clk
		.areset    (),                //        areset_conduit.export
		.locked    (),                //        locked_conduit.export
		.phasedone ()                 //     phasedone_conduit.export
	);

endmodule
