module Median_Filter (
    input  i_clk,
    input  i_rst_n
);
    
endmodule