module AudRecorder (
    input         i_rst_n, 
	input         i_clk,
	input         i_adclrck,
	input         i_en,
	input  [15:0] i_aud_adcdat,
	output [15:0] o_adc_data
);
    
endmodule
