module AudPlayer (
    input         i_rst_n,
	input         i_bclk,
	input         i_daclrck,
	input         i_en,
	input  [15:0] i_dac_data,
	output [15:0] o_aud_dacdat
);
    
endmodule
