module Corner_Finder (
    input  i_clk,
    input  i_rst_n
);
    
endmodule